library verilog;
use verilog.vl_types.all;
entity Index_Register_tb is
end Index_Register_tb;
