library verilog;
use verilog.vl_types.all;
entity girlanda_vlg_vec_tst is
end girlanda_vlg_vec_tst;
